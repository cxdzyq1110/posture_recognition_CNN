// megafunction wizard: %Shift register (RAM-based)%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSHIFT_TAPS 

// ============================================================
// File Name: line_buf_80pts_13lines.v
// Megafunction Name(s):
// 			ALTSHIFT_TAPS
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 14.0.0 Build 200 06/17/2014 SJ Full Version
// ************************************************************

//Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, the Altera Quartus II License Agreement,
//the Altera MegaCore Function License Agreement, or other 
//applicable license agreement, including, without limitation, 
//that your use is for the sole purpose of programming logic 
//devices manufactured by Altera and sold by Altera or its 
//authorized distributors.  Please refer to the applicable 
//agreement for further details.

module line_buf_80pts_13lines (
	aclr,
	clken,
	clock,
	shiftin,
	shiftout,
	taps0x,
	taps10x,
	taps11x,
	taps12x,
	taps1x,
	taps2x,
	taps3x,
	taps4x,
	taps5x,
	taps6x,
	taps7x,
	taps8x,
	taps9x);

	input	  aclr;
	input	  clken;
	input	  clock;
	input	[35:0]  shiftin;
	output	[35:0]  shiftout;
	output	[35:0]  taps0x;
	output	[35:0]  taps10x;
	output	[35:0]  taps11x;
	output	[35:0]  taps12x;
	output	[35:0]  taps1x;
	output	[35:0]  taps2x;
	output	[35:0]  taps3x;
	output	[35:0]  taps4x;
	output	[35:0]  taps5x;
	output	[35:0]  taps6x;
	output	[35:0]  taps7x;
	output	[35:0]  taps8x;
	output	[35:0]  taps9x;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  aclr;
	tri1	  clken;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACLR NUMERIC "1"
// Retrieval info: PRIVATE: CLKEN NUMERIC "1"
// Retrieval info: PRIVATE: GROUP_TAPS NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: NUMBER_OF_TAPS NUMERIC "13"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "1"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: TAP_DISTANCE NUMERIC "80"
// Retrieval info: PRIVATE: WIDTH NUMERIC "36"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: CONSTANT: LPM_HINT STRING "RAM_BLOCK_TYPE=M10K"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altshift_taps"
// Retrieval info: CONSTANT: NUMBER_OF_TAPS NUMERIC "13"
// Retrieval info: CONSTANT: TAP_DISTANCE NUMERIC "80"
// Retrieval info: CONSTANT: WIDTH NUMERIC "36"
// Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT VCC "aclr"
// Retrieval info: USED_PORT: clken 0 0 0 0 INPUT VCC "clken"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: shiftin 0 0 36 0 INPUT NODEFVAL "shiftin[35..0]"
// Retrieval info: USED_PORT: shiftout 0 0 36 0 OUTPUT NODEFVAL "shiftout[35..0]"
// Retrieval info: USED_PORT: taps0x 0 0 36 0 OUTPUT NODEFVAL "taps0x[35..0]"
// Retrieval info: USED_PORT: taps10x 0 0 36 0 OUTPUT NODEFVAL "taps10x[35..0]"
// Retrieval info: USED_PORT: taps11x 0 0 36 0 OUTPUT NODEFVAL "taps11x[35..0]"
// Retrieval info: USED_PORT: taps12x 0 0 36 0 OUTPUT NODEFVAL "taps12x[35..0]"
// Retrieval info: USED_PORT: taps1x 0 0 36 0 OUTPUT NODEFVAL "taps1x[35..0]"
// Retrieval info: USED_PORT: taps2x 0 0 36 0 OUTPUT NODEFVAL "taps2x[35..0]"
// Retrieval info: USED_PORT: taps3x 0 0 36 0 OUTPUT NODEFVAL "taps3x[35..0]"
// Retrieval info: USED_PORT: taps4x 0 0 36 0 OUTPUT NODEFVAL "taps4x[35..0]"
// Retrieval info: USED_PORT: taps5x 0 0 36 0 OUTPUT NODEFVAL "taps5x[35..0]"
// Retrieval info: USED_PORT: taps6x 0 0 36 0 OUTPUT NODEFVAL "taps6x[35..0]"
// Retrieval info: USED_PORT: taps7x 0 0 36 0 OUTPUT NODEFVAL "taps7x[35..0]"
// Retrieval info: USED_PORT: taps8x 0 0 36 0 OUTPUT NODEFVAL "taps8x[35..0]"
// Retrieval info: USED_PORT: taps9x 0 0 36 0 OUTPUT NODEFVAL "taps9x[35..0]"
// Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
// Retrieval info: CONNECT: @clken 0 0 0 0 clken 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @shiftin 0 0 36 0 shiftin 0 0 36 0
// Retrieval info: CONNECT: shiftout 0 0 36 0 @shiftout 0 0 36 0
// Retrieval info: CONNECT: taps0x 0 0 36 0 @taps 0 0 36 0
// Retrieval info: CONNECT: taps10x 0 0 36 0 @taps 0 0 36 360
// Retrieval info: CONNECT: taps11x 0 0 36 0 @taps 0 0 36 396
// Retrieval info: CONNECT: taps12x 0 0 36 0 @taps 0 0 36 432
// Retrieval info: CONNECT: taps1x 0 0 36 0 @taps 0 0 36 36
// Retrieval info: CONNECT: taps2x 0 0 36 0 @taps 0 0 36 72
// Retrieval info: CONNECT: taps3x 0 0 36 0 @taps 0 0 36 108
// Retrieval info: CONNECT: taps4x 0 0 36 0 @taps 0 0 36 144
// Retrieval info: CONNECT: taps5x 0 0 36 0 @taps 0 0 36 180
// Retrieval info: CONNECT: taps6x 0 0 36 0 @taps 0 0 36 216
// Retrieval info: CONNECT: taps7x 0 0 36 0 @taps 0 0 36 252
// Retrieval info: CONNECT: taps8x 0 0 36 0 @taps 0 0 36 288
// Retrieval info: CONNECT: taps9x 0 0 36 0 @taps 0 0 36 324
// Retrieval info: GEN_FILE: TYPE_NORMAL line_buf_80pts_13lines.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL line_buf_80pts_13lines.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL line_buf_80pts_13lines.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL line_buf_80pts_13lines.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL line_buf_80pts_13lines_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL line_buf_80pts_13lines_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
