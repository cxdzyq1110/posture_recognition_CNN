// soc_system.v

// Generated using ACDS version 14.0 200 at 2018.04.18.12:49:36

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        avalon_clk_clk,                       //                  avalon_clk.clk
		input  wire        avalon_reset_reset_n,                 //                avalon_reset.reset_n
		input  wire        avalon_clk_lw_clk,                    //               avalon_clk_lw.clk
		input  wire        avalon_reset_lw_reset_n,              //             avalon_reset_lw.reset_n
		output wire [14:0] memory_mem_a,                         //                      memory.mem_a
		output wire [2:0]  memory_mem_ba,                        //                            .mem_ba
		output wire        memory_mem_ck,                        //                            .mem_ck
		output wire        memory_mem_ck_n,                      //                            .mem_ck_n
		output wire        memory_mem_cke,                       //                            .mem_cke
		output wire        memory_mem_cs_n,                      //                            .mem_cs_n
		output wire        memory_mem_ras_n,                     //                            .mem_ras_n
		output wire        memory_mem_cas_n,                     //                            .mem_cas_n
		output wire        memory_mem_we_n,                      //                            .mem_we_n
		output wire        memory_mem_reset_n,                   //                            .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                        //                            .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                       //                            .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                     //                            .mem_dqs_n
		output wire        memory_mem_odt,                       //                            .mem_odt
		output wire [3:0]  memory_mem_dm,                        //                            .mem_dm
		input  wire        memory_oct_rzqin,                     //                            .oct_rzqin
		output wire        hps_io_hps_io_emac1_inst_TX_CLK,      //                      hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,        //                            .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,        //                            .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,        //                            .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,        //                            .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,        //                            .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,        //                            .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,         //                            .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL,      //                            .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL,      //                            .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK,      //                            .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,        //                            .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,        //                            .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,        //                            .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_sdio_inst_CMD,          //                            .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,           //                            .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,           //                            .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,          //                            .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,           //                            .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,           //                            .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,           //                            .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,           //                            .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,           //                            .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,           //                            .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,           //                            .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,           //                            .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,           //                            .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,           //                            .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,          //                            .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,          //                            .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,          //                            .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,          //                            .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,         //                            .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,        //                            .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,        //                            .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,         //                            .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,          //                            .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,          //                            .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,          //                            .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,          //                            .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,          //                            .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,          //                            .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,       //                            .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,       //                            .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO40,       //                            .hps_io_gpio_inst_GPIO40
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,       //                            .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,       //                            .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,       //                            .hps_io_gpio_inst_GPIO61
		input  wire        hps_0_f2h_cold_reset_req_reset_n,     //    hps_0_f2h_cold_reset_req.reset_n
		input  wire        hps_0_f2h_debug_reset_req_reset_n,    //   hps_0_f2h_debug_reset_req.reset_n
		input  wire [27:0] hps_0_f2h_stm_hw_events_stm_hwevents, //     hps_0_f2h_stm_hw_events.stm_hwevents
		input  wire        hps_0_f2h_warm_reset_req_reset_n,     //    hps_0_f2h_warm_reset_req.reset_n
		output wire        hps_0_h2f_reset_reset_n,              //             hps_0_h2f_reset.reset_n
		input  wire [29:0] avalon_f2s0_address,                  //                 avalon_f2s0.address
		input  wire [7:0]  avalon_f2s0_burstcount,               //                            .burstcount
		output wire        avalon_f2s0_waitrequest,              //                            .waitrequest
		output wire [31:0] avalon_f2s0_readdata,                 //                            .readdata
		output wire        avalon_f2s0_readdatavalid,            //                            .readdatavalid
		input  wire        avalon_f2s0_read,                     //                            .read
		input  wire [31:0] avalon_f2s0_writedata,                //                            .writedata
		input  wire [3:0]  avalon_f2s0_byteenable,               //                            .byteenable
		input  wire        avalon_f2s0_write,                    //                            .write
		output wire [7:0]  led_pio_external_connection_export,   // led_pio_external_connection.export
		input  wire [31:0] avalon_f2h_address,                   //                  avalon_f2h.address
		output wire        avalon_f2h_waitrequest,               //                            .waitrequest
		input  wire [3:0]  avalon_f2h_burstcount,                //                            .burstcount
		input  wire [3:0]  avalon_f2h_byteenable,                //                            .byteenable
		input  wire        avalon_f2h_beginbursttransfer,        //                            .beginbursttransfer
		input  wire        avalon_f2h_begintransfer,             //                            .begintransfer
		input  wire        avalon_f2h_read,                      //                            .read
		output wire [31:0] avalon_f2h_readdata,                  //                            .readdata
		output wire        avalon_f2h_readdatavalid,             //                            .readdatavalid
		input  wire        avalon_f2h_write,                     //                            .write
		input  wire [31:0] avalon_f2h_writedata,                 //                            .writedata
		output wire [21:0] avalon_h2f_address,                   //                  avalon_h2f.address
		output wire        avalon_h2f_write,                     //                            .write
		output wire        avalon_h2f_read,                      //                            .read
		input  wire [31:0] avalon_h2f_readdata,                  //                            .readdata
		output wire [31:0] avalon_h2f_writedata,                 //                            .writedata
		output wire        avalon_h2f_begintransfer,             //                            .begintransfer
		output wire        avalon_h2f_beginbursttransfer,        //                            .beginbursttransfer
		output wire [3:0]  avalon_h2f_burstcount,                //                            .burstcount
		output wire [3:0]  avalon_h2f_byteenable,                //                            .byteenable
		input  wire        avalon_h2f_readdatavalid,             //                            .readdatavalid
		input  wire        avalon_h2f_waitrequest,               //                            .waitrequest
		output wire [15:0] avalon_h2f_lw_address,                //               avalon_h2f_lw.address
		output wire        avalon_h2f_lw_write,                  //                            .write
		output wire        avalon_h2f_lw_read,                   //                            .read
		input  wire [31:0] avalon_h2f_lw_readdata,               //                            .readdata
		output wire [31:0] avalon_h2f_lw_writedata,              //                            .writedata
		output wire        avalon_h2f_lw_begintransfer,          //                            .begintransfer
		output wire        avalon_h2f_lw_beginbursttransfer,     //                            .beginbursttransfer
		output wire [3:0]  avalon_h2f_lw_burstcount,             //                            .burstcount
		output wire [3:0]  avalon_h2f_lw_byteenable,             //                            .byteenable
		input  wire        avalon_h2f_lw_readdatavalid,          //                            .readdatavalid
		input  wire        avalon_h2f_lw_waitrequest,            //                            .waitrequest
		input  wire [31:0] cnn_inst_info_export,                 //               cnn_inst_info.export
		input  wire [31:0] video_block_number_export,            //          video_block_number.export
		input  wire [29:0] avalon_f2s1_address,                  //                 avalon_f2s1.address
		input  wire [7:0]  avalon_f2s1_burstcount,               //                            .burstcount
		output wire        avalon_f2s1_waitrequest,              //                            .waitrequest
		output wire [31:0] avalon_f2s1_readdata,                 //                            .readdata
		output wire        avalon_f2s1_readdatavalid,            //                            .readdatavalid
		input  wire        avalon_f2s1_read,                     //                            .read
		input  wire [31:0] avalon_f2s1_writedata,                //                            .writedata
		input  wire [3:0]  avalon_f2s1_byteenable,               //                            .byteenable
		input  wire        avalon_f2s1_write,                    //                            .write
		output wire [7:0]  pd_bbox_frame_export,                 //               pd_bbox_frame.export
		output wire [11:0] pd_bbox_h2f_lw_address,               //              pd_bbox_h2f_lw.address
		output wire        pd_bbox_h2f_lw_write,                 //                            .write
		output wire        pd_bbox_h2f_lw_read,                  //                            .read
		input  wire [31:0] pd_bbox_h2f_lw_readdata,              //                            .readdata
		output wire [31:0] pd_bbox_h2f_lw_writedata,             //                            .writedata
		output wire        pd_bbox_h2f_lw_begintransfer,         //                            .begintransfer
		output wire        pd_bbox_h2f_lw_beginbursttransfer,    //                            .beginbursttransfer
		output wire [3:0]  pd_bbox_h2f_lw_burstcount,            //                            .burstcount
		output wire [3:0]  pd_bbox_h2f_lw_byteenable,            //                            .byteenable
		input  wire        pd_bbox_h2f_lw_readdatavalid,         //                            .readdatavalid
		input  wire        pd_bbox_h2f_lw_waitrequest,           //                            .waitrequest
		input  wire [29:0] avalon_f2s2_address,                  //                 avalon_f2s2.address
		input  wire [7:0]  avalon_f2s2_burstcount,               //                            .burstcount
		output wire        avalon_f2s2_waitrequest,              //                            .waitrequest
		output wire [31:0] avalon_f2s2_readdata,                 //                            .readdata
		output wire        avalon_f2s2_readdatavalid,            //                            .readdatavalid
		input  wire        avalon_f2s2_read,                     //                            .read
		input  wire [31:0] avalon_f2s2_writedata,                //                            .writedata
		input  wire [3:0]  avalon_f2s2_byteenable,               //                            .byteenable
		input  wire        avalon_f2s2_write                     //                            .write
	);

	wire          hps_0_h2f_lw_axi_master_awvalid;                                         // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                                          // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                                          // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                                         // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire          hps_0_h2f_lw_axi_master_arready;                                         // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                                            // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire          hps_0_h2f_lw_axi_master_rready;                                          // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire          hps_0_h2f_lw_axi_master_bready;                                          // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                                          // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                                          // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire          hps_0_h2f_lw_axi_master_arvalid;                                         // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                                          // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                                             // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                                           // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire          hps_0_h2f_lw_axi_master_awready;                                         // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                                            // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire          hps_0_h2f_lw_axi_master_bvalid;                                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                                             // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                                          // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                                         // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                                           // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_rvalid;                                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                                           // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_wready;                                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                                         // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                                          // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                                         // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                                           // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                                          // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                                             // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_wvalid;                                          // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire          hps_0_h2f_lw_axi_master_wlast;                                           // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire          hps_0_h2f_lw_axi_master_rlast;                                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire    [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;                    // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire   [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;                   // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [31:0] mm_interconnect_0_led_pio_s1_writedata;                                  // mm_interconnect_0:led_pio_s1_writedata -> led_pio:writedata
	wire    [1:0] mm_interconnect_0_led_pio_s1_address;                                    // mm_interconnect_0:led_pio_s1_address -> led_pio:address
	wire          mm_interconnect_0_led_pio_s1_chipselect;                                 // mm_interconnect_0:led_pio_s1_chipselect -> led_pio:chipselect
	wire          mm_interconnect_0_led_pio_s1_write;                                      // mm_interconnect_0:led_pio_s1_write -> led_pio:write_n
	wire   [31:0] mm_interconnect_0_led_pio_s1_readdata;                                   // led_pio:readdata -> mm_interconnect_0:led_pio_s1_readdata
	wire          mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_waitrequest;    // avalon_h2f_lw:uav_waitrequest -> mm_interconnect_0:avalon_h2f_lw_avalon_universal_slave_0_waitrequest
	wire    [3:0] mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_burstcount;     // mm_interconnect_0:avalon_h2f_lw_avalon_universal_slave_0_burstcount -> avalon_h2f_lw:uav_burstcount
	wire   [31:0] mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_writedata;      // mm_interconnect_0:avalon_h2f_lw_avalon_universal_slave_0_writedata -> avalon_h2f_lw:uav_writedata
	wire   [15:0] mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_address;        // mm_interconnect_0:avalon_h2f_lw_avalon_universal_slave_0_address -> avalon_h2f_lw:uav_address
	wire          mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_lock;           // mm_interconnect_0:avalon_h2f_lw_avalon_universal_slave_0_lock -> avalon_h2f_lw:uav_lock
	wire          mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_write;          // mm_interconnect_0:avalon_h2f_lw_avalon_universal_slave_0_write -> avalon_h2f_lw:uav_write
	wire          mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_read;           // mm_interconnect_0:avalon_h2f_lw_avalon_universal_slave_0_read -> avalon_h2f_lw:uav_read
	wire   [31:0] mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_readdata;       // avalon_h2f_lw:uav_readdata -> mm_interconnect_0:avalon_h2f_lw_avalon_universal_slave_0_readdata
	wire          mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_debugaccess;    // mm_interconnect_0:avalon_h2f_lw_avalon_universal_slave_0_debugaccess -> avalon_h2f_lw:uav_debugaccess
	wire          mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_readdatavalid;  // avalon_h2f_lw:uav_readdatavalid -> mm_interconnect_0:avalon_h2f_lw_avalon_universal_slave_0_readdatavalid
	wire    [3:0] mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_byteenable;     // mm_interconnect_0:avalon_h2f_lw_avalon_universal_slave_0_byteenable -> avalon_h2f_lw:uav_byteenable
	wire   [31:0] mm_interconnect_0_h2f_lw_ram_s1_writedata;                               // mm_interconnect_0:h2f_lw_ram_s1_writedata -> h2f_lw_ram:writedata
	wire    [1:0] mm_interconnect_0_h2f_lw_ram_s1_address;                                 // mm_interconnect_0:h2f_lw_ram_s1_address -> h2f_lw_ram:address
	wire          mm_interconnect_0_h2f_lw_ram_s1_chipselect;                              // mm_interconnect_0:h2f_lw_ram_s1_chipselect -> h2f_lw_ram:chipselect
	wire          mm_interconnect_0_h2f_lw_ram_s1_clken;                                   // mm_interconnect_0:h2f_lw_ram_s1_clken -> h2f_lw_ram:clken
	wire          mm_interconnect_0_h2f_lw_ram_s1_write;                                   // mm_interconnect_0:h2f_lw_ram_s1_write -> h2f_lw_ram:write
	wire   [31:0] mm_interconnect_0_h2f_lw_ram_s1_readdata;                                // h2f_lw_ram:readdata -> mm_interconnect_0:h2f_lw_ram_s1_readdata
	wire    [3:0] mm_interconnect_0_h2f_lw_ram_s1_byteenable;                              // mm_interconnect_0:h2f_lw_ram_s1_byteenable -> h2f_lw_ram:byteenable
	wire    [1:0] mm_interconnect_0_cnn_inst_info_s1_address;                              // mm_interconnect_0:cnn_inst_info_s1_address -> cnn_inst_info:address
	wire   [31:0] mm_interconnect_0_cnn_inst_info_s1_readdata;                             // cnn_inst_info:readdata -> mm_interconnect_0:cnn_inst_info_s1_readdata
	wire    [1:0] mm_interconnect_0_video_block_number_s1_address;                         // mm_interconnect_0:video_block_number_s1_address -> video_block_number:address
	wire   [31:0] mm_interconnect_0_video_block_number_s1_readdata;                        // video_block_number:readdata -> mm_interconnect_0:video_block_number_s1_readdata
	wire   [31:0] mm_interconnect_0_pd_bbox_frame_s1_writedata;                            // mm_interconnect_0:pd_bbox_frame_s1_writedata -> pd_bbox_frame:writedata
	wire    [1:0] mm_interconnect_0_pd_bbox_frame_s1_address;                              // mm_interconnect_0:pd_bbox_frame_s1_address -> pd_bbox_frame:address
	wire          mm_interconnect_0_pd_bbox_frame_s1_chipselect;                           // mm_interconnect_0:pd_bbox_frame_s1_chipselect -> pd_bbox_frame:chipselect
	wire          mm_interconnect_0_pd_bbox_frame_s1_write;                                // mm_interconnect_0:pd_bbox_frame_s1_write -> pd_bbox_frame:write_n
	wire   [31:0] mm_interconnect_0_pd_bbox_frame_s1_readdata;                             // pd_bbox_frame:readdata -> mm_interconnect_0:pd_bbox_frame_s1_readdata
	wire          mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_waitrequest;   // pd_bbox_h2f_lw:uav_waitrequest -> mm_interconnect_0:pd_bbox_h2f_lw_avalon_universal_slave_0_waitrequest
	wire    [3:0] mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_burstcount;    // mm_interconnect_0:pd_bbox_h2f_lw_avalon_universal_slave_0_burstcount -> pd_bbox_h2f_lw:uav_burstcount
	wire   [31:0] mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_writedata;     // mm_interconnect_0:pd_bbox_h2f_lw_avalon_universal_slave_0_writedata -> pd_bbox_h2f_lw:uav_writedata
	wire   [11:0] mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_address;       // mm_interconnect_0:pd_bbox_h2f_lw_avalon_universal_slave_0_address -> pd_bbox_h2f_lw:uav_address
	wire          mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_lock;          // mm_interconnect_0:pd_bbox_h2f_lw_avalon_universal_slave_0_lock -> pd_bbox_h2f_lw:uav_lock
	wire          mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_write;         // mm_interconnect_0:pd_bbox_h2f_lw_avalon_universal_slave_0_write -> pd_bbox_h2f_lw:uav_write
	wire          mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_read;          // mm_interconnect_0:pd_bbox_h2f_lw_avalon_universal_slave_0_read -> pd_bbox_h2f_lw:uav_read
	wire   [31:0] mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_readdata;      // pd_bbox_h2f_lw:uav_readdata -> mm_interconnect_0:pd_bbox_h2f_lw_avalon_universal_slave_0_readdata
	wire          mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_debugaccess;   // mm_interconnect_0:pd_bbox_h2f_lw_avalon_universal_slave_0_debugaccess -> pd_bbox_h2f_lw:uav_debugaccess
	wire          mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_readdatavalid; // pd_bbox_h2f_lw:uav_readdatavalid -> mm_interconnect_0:pd_bbox_h2f_lw_avalon_universal_slave_0_readdatavalid
	wire    [3:0] mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_byteenable;    // mm_interconnect_0:pd_bbox_h2f_lw_avalon_universal_slave_0_byteenable -> pd_bbox_h2f_lw:uav_byteenable
	wire          avalon_f2h_avalon_universal_master_0_waitrequest;                        // mm_interconnect_1:avalon_f2h_avalon_universal_master_0_waitrequest -> avalon_f2h:uav_waitrequest
	wire    [3:0] avalon_f2h_avalon_universal_master_0_burstcount;                         // avalon_f2h:uav_burstcount -> mm_interconnect_1:avalon_f2h_avalon_universal_master_0_burstcount
	wire   [31:0] avalon_f2h_avalon_universal_master_0_writedata;                          // avalon_f2h:uav_writedata -> mm_interconnect_1:avalon_f2h_avalon_universal_master_0_writedata
	wire   [31:0] avalon_f2h_avalon_universal_master_0_address;                            // avalon_f2h:uav_address -> mm_interconnect_1:avalon_f2h_avalon_universal_master_0_address
	wire          avalon_f2h_avalon_universal_master_0_lock;                               // avalon_f2h:uav_lock -> mm_interconnect_1:avalon_f2h_avalon_universal_master_0_lock
	wire          avalon_f2h_avalon_universal_master_0_write;                              // avalon_f2h:uav_write -> mm_interconnect_1:avalon_f2h_avalon_universal_master_0_write
	wire          avalon_f2h_avalon_universal_master_0_read;                               // avalon_f2h:uav_read -> mm_interconnect_1:avalon_f2h_avalon_universal_master_0_read
	wire   [31:0] avalon_f2h_avalon_universal_master_0_readdata;                           // mm_interconnect_1:avalon_f2h_avalon_universal_master_0_readdata -> avalon_f2h:uav_readdata
	wire          avalon_f2h_avalon_universal_master_0_debugaccess;                        // avalon_f2h:uav_debugaccess -> mm_interconnect_1:avalon_f2h_avalon_universal_master_0_debugaccess
	wire    [3:0] avalon_f2h_avalon_universal_master_0_byteenable;                         // avalon_f2h:uav_byteenable -> mm_interconnect_1:avalon_f2h_avalon_universal_master_0_byteenable
	wire          avalon_f2h_avalon_universal_master_0_readdatavalid;                      // mm_interconnect_1:avalon_f2h_avalon_universal_master_0_readdatavalid -> avalon_f2h:uav_readdatavalid
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_awvalid;                           // mm_interconnect_1:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire    [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_arsize;                            // mm_interconnect_1:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_arlock;                            // mm_interconnect_1:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire    [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_awcache;                           // mm_interconnect_1:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_arready;                           // hps_0:f2h_ARREADY -> mm_interconnect_1:hps_0_f2h_axi_slave_arready
	wire    [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_arid;                              // mm_interconnect_1:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_rready;                            // mm_interconnect_1:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_bready;                            // mm_interconnect_1:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire    [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_awsize;                            // mm_interconnect_1:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire    [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_awprot;                            // mm_interconnect_1:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_arvalid;                           // mm_interconnect_1:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire    [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_arprot;                            // mm_interconnect_1:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire    [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_bid;                               // hps_0:f2h_BID -> mm_interconnect_1:hps_0_f2h_axi_slave_bid
	wire    [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_arlen;                             // mm_interconnect_1:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_awready;                           // hps_0:f2h_AWREADY -> mm_interconnect_1:hps_0_f2h_axi_slave_awready
	wire    [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_awid;                              // mm_interconnect_1:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_bvalid;                            // hps_0:f2h_BVALID -> mm_interconnect_1:hps_0_f2h_axi_slave_bvalid
	wire    [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_wid;                               // mm_interconnect_1:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_awlock;                            // mm_interconnect_1:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_awburst;                           // mm_interconnect_1:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_bresp;                             // hps_0:f2h_BRESP -> mm_interconnect_1:hps_0_f2h_axi_slave_bresp
	wire    [4:0] mm_interconnect_1_hps_0_f2h_axi_slave_aruser;                            // mm_interconnect_1:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire    [4:0] mm_interconnect_1_hps_0_f2h_axi_slave_awuser;                            // mm_interconnect_1:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire    [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_wstrb;                             // mm_interconnect_1:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_rvalid;                            // hps_0:f2h_RVALID -> mm_interconnect_1:hps_0_f2h_axi_slave_rvalid
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_arburst;                           // mm_interconnect_1:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire   [31:0] mm_interconnect_1_hps_0_f2h_axi_slave_wdata;                             // mm_interconnect_1:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_wready;                            // hps_0:f2h_WREADY -> mm_interconnect_1:hps_0_f2h_axi_slave_wready
	wire   [31:0] mm_interconnect_1_hps_0_f2h_axi_slave_rdata;                             // hps_0:f2h_RDATA -> mm_interconnect_1:hps_0_f2h_axi_slave_rdata
	wire   [31:0] mm_interconnect_1_hps_0_f2h_axi_slave_araddr;                            // mm_interconnect_1:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire    [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_arcache;                           // mm_interconnect_1:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire    [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_awlen;                             // mm_interconnect_1:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire   [31:0] mm_interconnect_1_hps_0_f2h_axi_slave_awaddr;                            // mm_interconnect_1:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire    [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_rid;                               // hps_0:f2h_RID -> mm_interconnect_1:hps_0_f2h_axi_slave_rid
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_wvalid;                            // mm_interconnect_1:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_rresp;                             // hps_0:f2h_RRESP -> mm_interconnect_1:hps_0_f2h_axi_slave_rresp
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_wlast;                             // mm_interconnect_1:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_rlast;                             // hps_0:f2h_RLAST -> mm_interconnect_1:hps_0_f2h_axi_slave_rlast
	wire          hps_0_h2f_axi_master_awvalid;                                            // hps_0:h2f_AWVALID -> mm_interconnect_2:hps_0_h2f_axi_master_awvalid
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                             // hps_0:h2f_ARSIZE -> mm_interconnect_2:hps_0_h2f_axi_master_arsize
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                             // hps_0:h2f_ARLOCK -> mm_interconnect_2:hps_0_h2f_axi_master_arlock
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                            // hps_0:h2f_AWCACHE -> mm_interconnect_2:hps_0_h2f_axi_master_awcache
	wire          hps_0_h2f_axi_master_arready;                                            // mm_interconnect_2:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire   [11:0] hps_0_h2f_axi_master_arid;                                               // hps_0:h2f_ARID -> mm_interconnect_2:hps_0_h2f_axi_master_arid
	wire          hps_0_h2f_axi_master_rready;                                             // hps_0:h2f_RREADY -> mm_interconnect_2:hps_0_h2f_axi_master_rready
	wire          hps_0_h2f_axi_master_bready;                                             // hps_0:h2f_BREADY -> mm_interconnect_2:hps_0_h2f_axi_master_bready
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                             // hps_0:h2f_AWSIZE -> mm_interconnect_2:hps_0_h2f_axi_master_awsize
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                             // hps_0:h2f_AWPROT -> mm_interconnect_2:hps_0_h2f_axi_master_awprot
	wire          hps_0_h2f_axi_master_arvalid;                                            // hps_0:h2f_ARVALID -> mm_interconnect_2:hps_0_h2f_axi_master_arvalid
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                             // hps_0:h2f_ARPROT -> mm_interconnect_2:hps_0_h2f_axi_master_arprot
	wire   [11:0] hps_0_h2f_axi_master_bid;                                                // mm_interconnect_2:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                              // hps_0:h2f_ARLEN -> mm_interconnect_2:hps_0_h2f_axi_master_arlen
	wire          hps_0_h2f_axi_master_awready;                                            // mm_interconnect_2:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire   [11:0] hps_0_h2f_axi_master_awid;                                               // hps_0:h2f_AWID -> mm_interconnect_2:hps_0_h2f_axi_master_awid
	wire          hps_0_h2f_axi_master_bvalid;                                             // mm_interconnect_2:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire   [11:0] hps_0_h2f_axi_master_wid;                                                // hps_0:h2f_WID -> mm_interconnect_2:hps_0_h2f_axi_master_wid
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                             // hps_0:h2f_AWLOCK -> mm_interconnect_2:hps_0_h2f_axi_master_awlock
	wire    [1:0] hps_0_h2f_axi_master_awburst;                                            // hps_0:h2f_AWBURST -> mm_interconnect_2:hps_0_h2f_axi_master_awburst
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                              // mm_interconnect_2:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire    [3:0] hps_0_h2f_axi_master_wstrb;                                              // hps_0:h2f_WSTRB -> mm_interconnect_2:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_rvalid;                                             // mm_interconnect_2:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire   [31:0] hps_0_h2f_axi_master_wdata;                                              // hps_0:h2f_WDATA -> mm_interconnect_2:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_wready;                                             // mm_interconnect_2:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                            // hps_0:h2f_ARBURST -> mm_interconnect_2:hps_0_h2f_axi_master_arburst
	wire   [31:0] hps_0_h2f_axi_master_rdata;                                              // mm_interconnect_2:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                             // hps_0:h2f_ARADDR -> mm_interconnect_2:hps_0_h2f_axi_master_araddr
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                            // hps_0:h2f_ARCACHE -> mm_interconnect_2:hps_0_h2f_axi_master_arcache
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                              // hps_0:h2f_AWLEN -> mm_interconnect_2:hps_0_h2f_axi_master_awlen
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                             // hps_0:h2f_AWADDR -> mm_interconnect_2:hps_0_h2f_axi_master_awaddr
	wire   [11:0] hps_0_h2f_axi_master_rid;                                                // mm_interconnect_2:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_wvalid;                                             // hps_0:h2f_WVALID -> mm_interconnect_2:hps_0_h2f_axi_master_wvalid
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                              // mm_interconnect_2:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire          hps_0_h2f_axi_master_wlast;                                              // hps_0:h2f_WLAST -> mm_interconnect_2:hps_0_h2f_axi_master_wlast
	wire          hps_0_h2f_axi_master_rlast;                                              // mm_interconnect_2:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire          mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_waitrequest;       // avalon_h2f:uav_waitrequest -> mm_interconnect_2:avalon_h2f_avalon_universal_slave_0_waitrequest
	wire    [3:0] mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_burstcount;        // mm_interconnect_2:avalon_h2f_avalon_universal_slave_0_burstcount -> avalon_h2f:uav_burstcount
	wire   [31:0] mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_writedata;         // mm_interconnect_2:avalon_h2f_avalon_universal_slave_0_writedata -> avalon_h2f:uav_writedata
	wire   [21:0] mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_address;           // mm_interconnect_2:avalon_h2f_avalon_universal_slave_0_address -> avalon_h2f:uav_address
	wire          mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_lock;              // mm_interconnect_2:avalon_h2f_avalon_universal_slave_0_lock -> avalon_h2f:uav_lock
	wire          mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_write;             // mm_interconnect_2:avalon_h2f_avalon_universal_slave_0_write -> avalon_h2f:uav_write
	wire          mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_read;              // mm_interconnect_2:avalon_h2f_avalon_universal_slave_0_read -> avalon_h2f:uav_read
	wire   [31:0] mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_readdata;          // avalon_h2f:uav_readdata -> mm_interconnect_2:avalon_h2f_avalon_universal_slave_0_readdata
	wire          mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_debugaccess;       // mm_interconnect_2:avalon_h2f_avalon_universal_slave_0_debugaccess -> avalon_h2f:uav_debugaccess
	wire          mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_readdatavalid;     // avalon_h2f:uav_readdatavalid -> mm_interconnect_2:avalon_h2f_avalon_universal_slave_0_readdatavalid
	wire    [3:0] mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_byteenable;        // mm_interconnect_2:avalon_h2f_avalon_universal_slave_0_byteenable -> avalon_h2f:uav_byteenable
	wire  [127:0] mm_interconnect_2_h2f_ram_s1_writedata;                                  // mm_interconnect_2:h2f_ram_s1_writedata -> h2f_ram:writedata
	wire    [3:0] mm_interconnect_2_h2f_ram_s1_address;                                    // mm_interconnect_2:h2f_ram_s1_address -> h2f_ram:address
	wire          mm_interconnect_2_h2f_ram_s1_chipselect;                                 // mm_interconnect_2:h2f_ram_s1_chipselect -> h2f_ram:chipselect
	wire          mm_interconnect_2_h2f_ram_s1_clken;                                      // mm_interconnect_2:h2f_ram_s1_clken -> h2f_ram:clken
	wire          mm_interconnect_2_h2f_ram_s1_write;                                      // mm_interconnect_2:h2f_ram_s1_write -> h2f_ram:write
	wire  [127:0] mm_interconnect_2_h2f_ram_s1_readdata;                                   // h2f_ram:readdata -> mm_interconnect_2:h2f_ram_s1_readdata
	wire   [15:0] mm_interconnect_2_h2f_ram_s1_byteenable;                                 // mm_interconnect_2:h2f_ram_s1_byteenable -> h2f_ram:byteenable
	wire          rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [avalon_h2f:reset, avalon_h2f_lw:reset, cnn_inst_info:reset_n, h2f_lw_ram:reset, h2f_ram:reset, led_pio:reset_n, mm_interconnect_0:sysid_qsys_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:avalon_h2f_reset_reset_bridge_in_reset_reset, pd_bbox_frame:reset_n, pd_bbox_h2f_lw:reset, rst_translator:in_reset, sysid_qsys_0:reset_n, video_block_number:reset_n]
	wire          rst_controller_reset_out_reset_req;                                      // rst_controller:reset_req -> [h2f_lw_ram:reset_req, h2f_ram:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                                      // rst_controller_001:reset_out -> [avalon_f2h:reset, mm_interconnect_1:avalon_f2h_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_002_reset_out_reset;                                      // rst_controller_002:reset_out -> [mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_003_reset_out_reset;                                      // rst_controller_003:reset_out -> mm_interconnect_1:hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset

	soc_system_hps_0 #(
		.F2S_Width (1),
		.S2F_Width (1)
	) hps_0 (
		.f2h_cold_rst_req_n       (hps_0_f2h_cold_reset_req_reset_n),              //  f2h_cold_reset_req.reset_n
		.f2h_dbg_rst_req_n        (hps_0_f2h_debug_reset_req_reset_n),             // f2h_debug_reset_req.reset_n
		.f2h_warm_rst_req_n       (hps_0_f2h_warm_reset_req_reset_n),              //  f2h_warm_reset_req.reset_n
		.f2h_stm_hwevents         (hps_0_f2h_stm_hw_events_stm_hwevents),          //   f2h_stm_hw_events.stm_hwevents
		.mem_a                    (memory_mem_a),                                  //              memory.mem_a
		.mem_ba                   (memory_mem_ba),                                 //                    .mem_ba
		.mem_ck                   (memory_mem_ck),                                 //                    .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                               //                    .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                //                    .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                               //                    .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                              //                    .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                              //                    .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                               //                    .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                            //                    .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                 //                    .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                //                    .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                              //                    .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                //                    .mem_odt
		.mem_dm                   (memory_mem_dm),                                 //                    .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                              //                    .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),               //              hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),                 //                    .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),                 //                    .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),                 //                    .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),                 //                    .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),                 //                    .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),                 //                    .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),                  //                    .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),               //                    .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),               //                    .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),               //                    .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),                 //                    .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),                 //                    .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),                 //                    .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),                   //                    .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),                    //                    .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),                    //                    .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),                   //                    .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),                    //                    .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),                    //                    .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),                    //                    .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),                    //                    .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),                    //                    .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),                    //                    .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),                    //                    .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),                    //                    .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),                    //                    .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),                    //                    .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),                   //                    .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),                   //                    .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),                   //                    .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),                   //                    .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),                  //                    .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),                 //                    .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),                 //                    .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),                  //                    .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),                   //                    .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),                   //                    .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),                   //                    .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),                   //                    .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),                   //                    .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),                   //                    .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),                //                    .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),                //                    .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),                //                    .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),                //                    .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),                //                    .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),                //                    .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),                       //           h2f_reset.reset_n
		.f2h_sdram0_clk           (avalon_clk_clk),                                //    f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (avalon_f2s0_address),                           //     f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (avalon_f2s0_burstcount),                        //                    .burstcount
		.f2h_sdram0_WAITREQUEST   (avalon_f2s0_waitrequest),                       //                    .waitrequest
		.f2h_sdram0_READDATA      (avalon_f2s0_readdata),                          //                    .readdata
		.f2h_sdram0_READDATAVALID (avalon_f2s0_readdatavalid),                     //                    .readdatavalid
		.f2h_sdram0_READ          (avalon_f2s0_read),                              //                    .read
		.f2h_sdram0_WRITEDATA     (avalon_f2s0_writedata),                         //                    .writedata
		.f2h_sdram0_BYTEENABLE    (avalon_f2s0_byteenable),                        //                    .byteenable
		.f2h_sdram0_WRITE         (avalon_f2s0_write),                             //                    .write
		.f2h_sdram1_clk           (avalon_clk_clk),                                //    f2h_sdram1_clock.clk
		.f2h_sdram1_ADDRESS       (avalon_f2s1_address),                           //     f2h_sdram1_data.address
		.f2h_sdram1_BURSTCOUNT    (avalon_f2s1_burstcount),                        //                    .burstcount
		.f2h_sdram1_WAITREQUEST   (avalon_f2s1_waitrequest),                       //                    .waitrequest
		.f2h_sdram1_READDATA      (avalon_f2s1_readdata),                          //                    .readdata
		.f2h_sdram1_READDATAVALID (avalon_f2s1_readdatavalid),                     //                    .readdatavalid
		.f2h_sdram1_READ          (avalon_f2s1_read),                              //                    .read
		.f2h_sdram1_WRITEDATA     (avalon_f2s1_writedata),                         //                    .writedata
		.f2h_sdram1_BYTEENABLE    (avalon_f2s1_byteenable),                        //                    .byteenable
		.f2h_sdram1_WRITE         (avalon_f2s1_write),                             //                    .write
		.f2h_sdram2_clk           (avalon_clk_clk),                                //    f2h_sdram2_clock.clk
		.f2h_sdram2_ADDRESS       (avalon_f2s2_address),                           //     f2h_sdram2_data.address
		.f2h_sdram2_BURSTCOUNT    (avalon_f2s2_burstcount),                        //                    .burstcount
		.f2h_sdram2_WAITREQUEST   (avalon_f2s2_waitrequest),                       //                    .waitrequest
		.f2h_sdram2_READDATA      (avalon_f2s2_readdata),                          //                    .readdata
		.f2h_sdram2_READDATAVALID (avalon_f2s2_readdatavalid),                     //                    .readdatavalid
		.f2h_sdram2_READ          (avalon_f2s2_read),                              //                    .read
		.f2h_sdram2_WRITEDATA     (avalon_f2s2_writedata),                         //                    .writedata
		.f2h_sdram2_BYTEENABLE    (avalon_f2s2_byteenable),                        //                    .byteenable
		.f2h_sdram2_WRITE         (avalon_f2s2_write),                             //                    .write
		.h2f_axi_clk              (avalon_clk_lw_clk),                             //       h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),                     //      h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),                   //                    .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),                    //                    .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),                   //                    .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),                  //                    .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),                   //                    .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),                  //                    .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),                   //                    .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),                  //                    .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),                  //                    .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),                      //                    .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),                    //                    .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),                    //                    .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),                    //                    .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),                   //                    .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),                   //                    .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),                      //                    .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),                    //                    .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),                   //                    .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),                   //                    .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),                     //                    .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),                   //                    .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),                    //                    .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),                   //                    .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),                  //                    .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),                   //                    .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),                  //                    .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),                   //                    .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),                  //                    .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),                  //                    .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),                      //                    .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),                    //                    .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),                    //                    .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),                    //                    .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),                   //                    .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),                   //                    .rready
		.f2h_axi_clk              (avalon_clk_clk),                                //       f2h_axi_clock.clk
		.f2h_AWID                 (mm_interconnect_1_hps_0_f2h_axi_slave_awid),    //       f2h_axi_slave.awid
		.f2h_AWADDR               (mm_interconnect_1_hps_0_f2h_axi_slave_awaddr),  //                    .awaddr
		.f2h_AWLEN                (mm_interconnect_1_hps_0_f2h_axi_slave_awlen),   //                    .awlen
		.f2h_AWSIZE               (mm_interconnect_1_hps_0_f2h_axi_slave_awsize),  //                    .awsize
		.f2h_AWBURST              (mm_interconnect_1_hps_0_f2h_axi_slave_awburst), //                    .awburst
		.f2h_AWLOCK               (mm_interconnect_1_hps_0_f2h_axi_slave_awlock),  //                    .awlock
		.f2h_AWCACHE              (mm_interconnect_1_hps_0_f2h_axi_slave_awcache), //                    .awcache
		.f2h_AWPROT               (mm_interconnect_1_hps_0_f2h_axi_slave_awprot),  //                    .awprot
		.f2h_AWVALID              (mm_interconnect_1_hps_0_f2h_axi_slave_awvalid), //                    .awvalid
		.f2h_AWREADY              (mm_interconnect_1_hps_0_f2h_axi_slave_awready), //                    .awready
		.f2h_AWUSER               (mm_interconnect_1_hps_0_f2h_axi_slave_awuser),  //                    .awuser
		.f2h_WID                  (mm_interconnect_1_hps_0_f2h_axi_slave_wid),     //                    .wid
		.f2h_WDATA                (mm_interconnect_1_hps_0_f2h_axi_slave_wdata),   //                    .wdata
		.f2h_WSTRB                (mm_interconnect_1_hps_0_f2h_axi_slave_wstrb),   //                    .wstrb
		.f2h_WLAST                (mm_interconnect_1_hps_0_f2h_axi_slave_wlast),   //                    .wlast
		.f2h_WVALID               (mm_interconnect_1_hps_0_f2h_axi_slave_wvalid),  //                    .wvalid
		.f2h_WREADY               (mm_interconnect_1_hps_0_f2h_axi_slave_wready),  //                    .wready
		.f2h_BID                  (mm_interconnect_1_hps_0_f2h_axi_slave_bid),     //                    .bid
		.f2h_BRESP                (mm_interconnect_1_hps_0_f2h_axi_slave_bresp),   //                    .bresp
		.f2h_BVALID               (mm_interconnect_1_hps_0_f2h_axi_slave_bvalid),  //                    .bvalid
		.f2h_BREADY               (mm_interconnect_1_hps_0_f2h_axi_slave_bready),  //                    .bready
		.f2h_ARID                 (mm_interconnect_1_hps_0_f2h_axi_slave_arid),    //                    .arid
		.f2h_ARADDR               (mm_interconnect_1_hps_0_f2h_axi_slave_araddr),  //                    .araddr
		.f2h_ARLEN                (mm_interconnect_1_hps_0_f2h_axi_slave_arlen),   //                    .arlen
		.f2h_ARSIZE               (mm_interconnect_1_hps_0_f2h_axi_slave_arsize),  //                    .arsize
		.f2h_ARBURST              (mm_interconnect_1_hps_0_f2h_axi_slave_arburst), //                    .arburst
		.f2h_ARLOCK               (mm_interconnect_1_hps_0_f2h_axi_slave_arlock),  //                    .arlock
		.f2h_ARCACHE              (mm_interconnect_1_hps_0_f2h_axi_slave_arcache), //                    .arcache
		.f2h_ARPROT               (mm_interconnect_1_hps_0_f2h_axi_slave_arprot),  //                    .arprot
		.f2h_ARVALID              (mm_interconnect_1_hps_0_f2h_axi_slave_arvalid), //                    .arvalid
		.f2h_ARREADY              (mm_interconnect_1_hps_0_f2h_axi_slave_arready), //                    .arready
		.f2h_ARUSER               (mm_interconnect_1_hps_0_f2h_axi_slave_aruser),  //                    .aruser
		.f2h_RID                  (mm_interconnect_1_hps_0_f2h_axi_slave_rid),     //                    .rid
		.f2h_RDATA                (mm_interconnect_1_hps_0_f2h_axi_slave_rdata),   //                    .rdata
		.f2h_RRESP                (mm_interconnect_1_hps_0_f2h_axi_slave_rresp),   //                    .rresp
		.f2h_RLAST                (mm_interconnect_1_hps_0_f2h_axi_slave_rlast),   //                    .rlast
		.f2h_RVALID               (mm_interconnect_1_hps_0_f2h_axi_slave_rvalid),  //                    .rvalid
		.f2h_RREADY               (mm_interconnect_1_hps_0_f2h_axi_slave_rready),  //                    .rready
		.h2f_lw_axi_clk           (avalon_clk_lw_clk),                             //    h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                  //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                //                    .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                 //                    .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                //                    .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),               //                    .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                //                    .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),               //                    .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                //                    .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),               //                    .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),               //                    .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                   //                    .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                 //                    .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                 //                    .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                 //                    .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                //                    .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                //                    .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                   //                    .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                 //                    .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                //                    .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                //                    .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                  //                    .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                //                    .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                 //                    .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                //                    .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),               //                    .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                //                    .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),               //                    .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                //                    .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),               //                    .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),               //                    .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                   //                    .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                 //                    .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                 //                    .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                 //                    .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                //                    .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready)                 //                    .rready
	);

	soc_system_sysid_qsys_0 sysid_qsys_0 (
		.clock    (avalon_clk_lw_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	soc_system_led_pio led_pio (
		.clk        (avalon_clk_lw_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_external_connection_export)       // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (4),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (4),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (1),
		.USE_BEGINTRANSFER           (1),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (0),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) avalon_f2h (
		.clk                      (avalon_clk_clk),                                     //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                 //                     reset.reset
		.uav_address              (avalon_f2h_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (avalon_f2h_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (avalon_f2h_avalon_universal_master_0_read),          //                          .read
		.uav_write                (avalon_f2h_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (avalon_f2h_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (avalon_f2h_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (avalon_f2h_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (avalon_f2h_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (avalon_f2h_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (avalon_f2h_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (avalon_f2h_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (avalon_f2h_address),                                 //      avalon_anti_master_0.address
		.av_waitrequest           (avalon_f2h_waitrequest),                             //                          .waitrequest
		.av_burstcount            (avalon_f2h_burstcount),                              //                          .burstcount
		.av_byteenable            (avalon_f2h_byteenable),                              //                          .byteenable
		.av_beginbursttransfer    (avalon_f2h_beginbursttransfer),                      //                          .beginbursttransfer
		.av_begintransfer         (avalon_f2h_begintransfer),                           //                          .begintransfer
		.av_read                  (avalon_f2h_read),                                    //                          .read
		.av_readdata              (avalon_f2h_readdata),                                //                          .readdata
		.av_readdatavalid         (avalon_f2h_readdatavalid),                           //                          .readdatavalid
		.av_write                 (avalon_f2h_write),                                   //                          .write
		.av_writedata             (avalon_f2h_writedata),                               //                          .writedata
		.av_chipselect            (1'b0),                                               //               (terminated)
		.av_lock                  (1'b0),                                               //               (terminated)
		.av_debugaccess           (1'b0),                                               //               (terminated)
		.uav_clken                (),                                                   //               (terminated)
		.av_clken                 (1'b1),                                               //               (terminated)
		.uav_response             (2'b00),                                              //               (terminated)
		.av_response              (),                                                   //               (terminated)
		.uav_writeresponserequest (),                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                               //               (terminated)
		.av_writeresponsevalid    ()                                                    //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (22),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (4),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (22),
		.UAV_BURSTCOUNT_W               (4),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) avalon_h2f (
		.clk                      (avalon_clk_lw_clk),                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                      //                    reset.reset
		.uav_address              (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_burstcount),    //                         .burstcount
		.uav_read                 (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_read),          //                         .read
		.uav_write                (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_write),         //                         .write
		.uav_waitrequest          (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_byteenable),    //                         .byteenable
		.uav_readdata             (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_readdata),      //                         .readdata
		.uav_writedata            (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_writedata),     //                         .writedata
		.uav_lock                 (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_lock),          //                         .lock
		.uav_debugaccess          (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_debugaccess),   //                         .debugaccess
		.av_address               (avalon_h2f_address),                                                  //      avalon_anti_slave_0.address
		.av_write                 (avalon_h2f_write),                                                    //                         .write
		.av_read                  (avalon_h2f_read),                                                     //                         .read
		.av_readdata              (avalon_h2f_readdata),                                                 //                         .readdata
		.av_writedata             (avalon_h2f_writedata),                                                //                         .writedata
		.av_begintransfer         (avalon_h2f_begintransfer),                                            //                         .begintransfer
		.av_beginbursttransfer    (avalon_h2f_beginbursttransfer),                                       //                         .beginbursttransfer
		.av_burstcount            (avalon_h2f_burstcount),                                               //                         .burstcount
		.av_byteenable            (avalon_h2f_byteenable),                                               //                         .byteenable
		.av_readdatavalid         (avalon_h2f_readdatavalid),                                            //                         .readdatavalid
		.av_waitrequest           (avalon_h2f_waitrequest),                                              //                         .waitrequest
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_chipselect            (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (16),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (4),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (16),
		.UAV_BURSTCOUNT_W               (4),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) avalon_h2f_lw (
		.clk                      (avalon_clk_lw_clk),                                                      //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address              (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_burstcount),    //                         .burstcount
		.uav_read                 (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_read),          //                         .read
		.uav_write                (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_write),         //                         .write
		.uav_waitrequest          (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_byteenable),    //                         .byteenable
		.uav_readdata             (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_readdata),      //                         .readdata
		.uav_writedata            (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_writedata),     //                         .writedata
		.uav_lock                 (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_lock),          //                         .lock
		.uav_debugaccess          (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_debugaccess),   //                         .debugaccess
		.av_address               (avalon_h2f_lw_address),                                                  //      avalon_anti_slave_0.address
		.av_write                 (avalon_h2f_lw_write),                                                    //                         .write
		.av_read                  (avalon_h2f_lw_read),                                                     //                         .read
		.av_readdata              (avalon_h2f_lw_readdata),                                                 //                         .readdata
		.av_writedata             (avalon_h2f_lw_writedata),                                                //                         .writedata
		.av_begintransfer         (avalon_h2f_lw_begintransfer),                                            //                         .begintransfer
		.av_beginbursttransfer    (avalon_h2f_lw_beginbursttransfer),                                       //                         .beginbursttransfer
		.av_burstcount            (avalon_h2f_lw_burstcount),                                               //                         .burstcount
		.av_byteenable            (avalon_h2f_lw_byteenable),                                               //                         .byteenable
		.av_readdatavalid         (avalon_h2f_lw_readdatavalid),                                            //                         .readdatavalid
		.av_waitrequest           (avalon_h2f_lw_waitrequest),                                              //                         .waitrequest
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	soc_system_h2f_ram h2f_ram (
		.clk        (avalon_clk_lw_clk),                       //   clk1.clk
		.address    (mm_interconnect_2_h2f_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_2_h2f_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_2_h2f_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_2_h2f_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_2_h2f_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_2_h2f_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_2_h2f_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)       //       .reset_req
	);

	soc_system_h2f_lw_ram h2f_lw_ram (
		.clk        (avalon_clk_lw_clk),                          //   clk1.clk
		.address    (mm_interconnect_0_h2f_lw_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_h2f_lw_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_h2f_lw_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_h2f_lw_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_h2f_lw_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_h2f_lw_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_h2f_lw_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)          //       .reset_req
	);

	soc_system_cnn_inst_info cnn_inst_info (
		.clk      (avalon_clk_lw_clk),                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_cnn_inst_info_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_cnn_inst_info_s1_readdata), //                    .readdata
		.in_port  (cnn_inst_info_export)                         // external_connection.export
	);

	soc_system_cnn_inst_info video_block_number (
		.clk      (avalon_clk_lw_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address  (mm_interconnect_0_video_block_number_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_video_block_number_s1_readdata), //                    .readdata
		.in_port  (video_block_number_export)                         // external_connection.export
	);

	soc_system_led_pio pd_bbox_frame (
		.clk        (avalon_clk_lw_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pd_bbox_frame_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pd_bbox_frame_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pd_bbox_frame_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pd_bbox_frame_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pd_bbox_frame_s1_readdata),   //                    .readdata
		.out_port   (pd_bbox_frame_export)                           // external_connection.export
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (12),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (4),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (12),
		.UAV_BURSTCOUNT_W               (4),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pd_bbox_h2f_lw (
		.clk                      (avalon_clk_lw_clk),                                                       //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address              (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_burstcount),    //                         .burstcount
		.uav_read                 (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_read),          //                         .read
		.uav_write                (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_write),         //                         .write
		.uav_waitrequest          (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_byteenable),    //                         .byteenable
		.uav_readdata             (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_readdata),      //                         .readdata
		.uav_writedata            (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_writedata),     //                         .writedata
		.uav_lock                 (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_lock),          //                         .lock
		.uav_debugaccess          (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_debugaccess),   //                         .debugaccess
		.av_address               (pd_bbox_h2f_lw_address),                                                  //      avalon_anti_slave_0.address
		.av_write                 (pd_bbox_h2f_lw_write),                                                    //                         .write
		.av_read                  (pd_bbox_h2f_lw_read),                                                     //                         .read
		.av_readdata              (pd_bbox_h2f_lw_readdata),                                                 //                         .readdata
		.av_writedata             (pd_bbox_h2f_lw_writedata),                                                //                         .writedata
		.av_begintransfer         (pd_bbox_h2f_lw_begintransfer),                                            //                         .begintransfer
		.av_beginbursttransfer    (pd_bbox_h2f_lw_beginbursttransfer),                                       //                         .beginbursttransfer
		.av_burstcount            (pd_bbox_h2f_lw_burstcount),                                               //                         .burstcount
		.av_byteenable            (pd_bbox_h2f_lw_byteenable),                                               //                         .byteenable
		.av_readdatavalid         (pd_bbox_h2f_lw_readdatavalid),                                            //                         .readdatavalid
		.av_waitrequest           (pd_bbox_h2f_lw_waitrequest),                                              //                         .waitrequest
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_chipselect            (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                                            //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                                          //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                                           //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                                          //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                                         //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                                          //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                                         //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                                          //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                                         //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                                         //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                                             //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                                           //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                                           //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                                           //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                                          //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                                          //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                                             //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                                           //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                                          //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                                          //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                                            //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                                          //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                                           //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                                          //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                                         //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                                          //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                                         //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                                          //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                                         //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                                         //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                                             //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                                           //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                                           //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                                           //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                                          //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                                          //                                                              .rready
		.clk_1_clk_clk                                                       (avalon_clk_lw_clk),                                                       //                                                     clk_1_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                      // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.sysid_qsys_0_reset_reset_bridge_in_reset_reset                      (rst_controller_reset_out_reset),                                          //                      sysid_qsys_0_reset_reset_bridge_in_reset.reset
		.avalon_h2f_lw_avalon_universal_slave_0_address                      (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_address),        //                        avalon_h2f_lw_avalon_universal_slave_0.address
		.avalon_h2f_lw_avalon_universal_slave_0_write                        (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_write),          //                                                              .write
		.avalon_h2f_lw_avalon_universal_slave_0_read                         (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_read),           //                                                              .read
		.avalon_h2f_lw_avalon_universal_slave_0_readdata                     (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_readdata),       //                                                              .readdata
		.avalon_h2f_lw_avalon_universal_slave_0_writedata                    (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_writedata),      //                                                              .writedata
		.avalon_h2f_lw_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_burstcount),     //                                                              .burstcount
		.avalon_h2f_lw_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_byteenable),     //                                                              .byteenable
		.avalon_h2f_lw_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_readdatavalid),  //                                                              .readdatavalid
		.avalon_h2f_lw_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_waitrequest),    //                                                              .waitrequest
		.avalon_h2f_lw_avalon_universal_slave_0_lock                         (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_lock),           //                                                              .lock
		.avalon_h2f_lw_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_avalon_h2f_lw_avalon_universal_slave_0_debugaccess),    //                                                              .debugaccess
		.cnn_inst_info_s1_address                                            (mm_interconnect_0_cnn_inst_info_s1_address),                              //                                              cnn_inst_info_s1.address
		.cnn_inst_info_s1_readdata                                           (mm_interconnect_0_cnn_inst_info_s1_readdata),                             //                                                              .readdata
		.h2f_lw_ram_s1_address                                               (mm_interconnect_0_h2f_lw_ram_s1_address),                                 //                                                 h2f_lw_ram_s1.address
		.h2f_lw_ram_s1_write                                                 (mm_interconnect_0_h2f_lw_ram_s1_write),                                   //                                                              .write
		.h2f_lw_ram_s1_readdata                                              (mm_interconnect_0_h2f_lw_ram_s1_readdata),                                //                                                              .readdata
		.h2f_lw_ram_s1_writedata                                             (mm_interconnect_0_h2f_lw_ram_s1_writedata),                               //                                                              .writedata
		.h2f_lw_ram_s1_byteenable                                            (mm_interconnect_0_h2f_lw_ram_s1_byteenable),                              //                                                              .byteenable
		.h2f_lw_ram_s1_chipselect                                            (mm_interconnect_0_h2f_lw_ram_s1_chipselect),                              //                                                              .chipselect
		.h2f_lw_ram_s1_clken                                                 (mm_interconnect_0_h2f_lw_ram_s1_clken),                                   //                                                              .clken
		.led_pio_s1_address                                                  (mm_interconnect_0_led_pio_s1_address),                                    //                                                    led_pio_s1.address
		.led_pio_s1_write                                                    (mm_interconnect_0_led_pio_s1_write),                                      //                                                              .write
		.led_pio_s1_readdata                                                 (mm_interconnect_0_led_pio_s1_readdata),                                   //                                                              .readdata
		.led_pio_s1_writedata                                                (mm_interconnect_0_led_pio_s1_writedata),                                  //                                                              .writedata
		.led_pio_s1_chipselect                                               (mm_interconnect_0_led_pio_s1_chipselect),                                 //                                                              .chipselect
		.pd_bbox_frame_s1_address                                            (mm_interconnect_0_pd_bbox_frame_s1_address),                              //                                              pd_bbox_frame_s1.address
		.pd_bbox_frame_s1_write                                              (mm_interconnect_0_pd_bbox_frame_s1_write),                                //                                                              .write
		.pd_bbox_frame_s1_readdata                                           (mm_interconnect_0_pd_bbox_frame_s1_readdata),                             //                                                              .readdata
		.pd_bbox_frame_s1_writedata                                          (mm_interconnect_0_pd_bbox_frame_s1_writedata),                            //                                                              .writedata
		.pd_bbox_frame_s1_chipselect                                         (mm_interconnect_0_pd_bbox_frame_s1_chipselect),                           //                                                              .chipselect
		.pd_bbox_h2f_lw_avalon_universal_slave_0_address                     (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_address),       //                       pd_bbox_h2f_lw_avalon_universal_slave_0.address
		.pd_bbox_h2f_lw_avalon_universal_slave_0_write                       (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_write),         //                                                              .write
		.pd_bbox_h2f_lw_avalon_universal_slave_0_read                        (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_read),          //                                                              .read
		.pd_bbox_h2f_lw_avalon_universal_slave_0_readdata                    (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_readdata),      //                                                              .readdata
		.pd_bbox_h2f_lw_avalon_universal_slave_0_writedata                   (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_writedata),     //                                                              .writedata
		.pd_bbox_h2f_lw_avalon_universal_slave_0_burstcount                  (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_burstcount),    //                                                              .burstcount
		.pd_bbox_h2f_lw_avalon_universal_slave_0_byteenable                  (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_byteenable),    //                                                              .byteenable
		.pd_bbox_h2f_lw_avalon_universal_slave_0_readdatavalid               (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_readdatavalid), //                                                              .readdatavalid
		.pd_bbox_h2f_lw_avalon_universal_slave_0_waitrequest                 (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_waitrequest),   //                                                              .waitrequest
		.pd_bbox_h2f_lw_avalon_universal_slave_0_lock                        (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_lock),          //                                                              .lock
		.pd_bbox_h2f_lw_avalon_universal_slave_0_debugaccess                 (mm_interconnect_0_pd_bbox_h2f_lw_avalon_universal_slave_0_debugaccess),   //                                                              .debugaccess
		.sysid_qsys_0_control_slave_address                                  (mm_interconnect_0_sysid_qsys_0_control_slave_address),                    //                                    sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                                 (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),                   //                                                              .readdata
		.video_block_number_s1_address                                       (mm_interconnect_0_video_block_number_s1_address),                         //                                         video_block_number_s1.address
		.video_block_number_s1_readdata                                      (mm_interconnect_0_video_block_number_s1_readdata)                         //                                                              .readdata
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_f2h_axi_slave_awid                                         (mm_interconnect_1_hps_0_f2h_axi_slave_awid),         //                                        hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                                       (mm_interconnect_1_hps_0_f2h_axi_slave_awaddr),       //                                                           .awaddr
		.hps_0_f2h_axi_slave_awlen                                        (mm_interconnect_1_hps_0_f2h_axi_slave_awlen),        //                                                           .awlen
		.hps_0_f2h_axi_slave_awsize                                       (mm_interconnect_1_hps_0_f2h_axi_slave_awsize),       //                                                           .awsize
		.hps_0_f2h_axi_slave_awburst                                      (mm_interconnect_1_hps_0_f2h_axi_slave_awburst),      //                                                           .awburst
		.hps_0_f2h_axi_slave_awlock                                       (mm_interconnect_1_hps_0_f2h_axi_slave_awlock),       //                                                           .awlock
		.hps_0_f2h_axi_slave_awcache                                      (mm_interconnect_1_hps_0_f2h_axi_slave_awcache),      //                                                           .awcache
		.hps_0_f2h_axi_slave_awprot                                       (mm_interconnect_1_hps_0_f2h_axi_slave_awprot),       //                                                           .awprot
		.hps_0_f2h_axi_slave_awuser                                       (mm_interconnect_1_hps_0_f2h_axi_slave_awuser),       //                                                           .awuser
		.hps_0_f2h_axi_slave_awvalid                                      (mm_interconnect_1_hps_0_f2h_axi_slave_awvalid),      //                                                           .awvalid
		.hps_0_f2h_axi_slave_awready                                      (mm_interconnect_1_hps_0_f2h_axi_slave_awready),      //                                                           .awready
		.hps_0_f2h_axi_slave_wid                                          (mm_interconnect_1_hps_0_f2h_axi_slave_wid),          //                                                           .wid
		.hps_0_f2h_axi_slave_wdata                                        (mm_interconnect_1_hps_0_f2h_axi_slave_wdata),        //                                                           .wdata
		.hps_0_f2h_axi_slave_wstrb                                        (mm_interconnect_1_hps_0_f2h_axi_slave_wstrb),        //                                                           .wstrb
		.hps_0_f2h_axi_slave_wlast                                        (mm_interconnect_1_hps_0_f2h_axi_slave_wlast),        //                                                           .wlast
		.hps_0_f2h_axi_slave_wvalid                                       (mm_interconnect_1_hps_0_f2h_axi_slave_wvalid),       //                                                           .wvalid
		.hps_0_f2h_axi_slave_wready                                       (mm_interconnect_1_hps_0_f2h_axi_slave_wready),       //                                                           .wready
		.hps_0_f2h_axi_slave_bid                                          (mm_interconnect_1_hps_0_f2h_axi_slave_bid),          //                                                           .bid
		.hps_0_f2h_axi_slave_bresp                                        (mm_interconnect_1_hps_0_f2h_axi_slave_bresp),        //                                                           .bresp
		.hps_0_f2h_axi_slave_bvalid                                       (mm_interconnect_1_hps_0_f2h_axi_slave_bvalid),       //                                                           .bvalid
		.hps_0_f2h_axi_slave_bready                                       (mm_interconnect_1_hps_0_f2h_axi_slave_bready),       //                                                           .bready
		.hps_0_f2h_axi_slave_arid                                         (mm_interconnect_1_hps_0_f2h_axi_slave_arid),         //                                                           .arid
		.hps_0_f2h_axi_slave_araddr                                       (mm_interconnect_1_hps_0_f2h_axi_slave_araddr),       //                                                           .araddr
		.hps_0_f2h_axi_slave_arlen                                        (mm_interconnect_1_hps_0_f2h_axi_slave_arlen),        //                                                           .arlen
		.hps_0_f2h_axi_slave_arsize                                       (mm_interconnect_1_hps_0_f2h_axi_slave_arsize),       //                                                           .arsize
		.hps_0_f2h_axi_slave_arburst                                      (mm_interconnect_1_hps_0_f2h_axi_slave_arburst),      //                                                           .arburst
		.hps_0_f2h_axi_slave_arlock                                       (mm_interconnect_1_hps_0_f2h_axi_slave_arlock),       //                                                           .arlock
		.hps_0_f2h_axi_slave_arcache                                      (mm_interconnect_1_hps_0_f2h_axi_slave_arcache),      //                                                           .arcache
		.hps_0_f2h_axi_slave_arprot                                       (mm_interconnect_1_hps_0_f2h_axi_slave_arprot),       //                                                           .arprot
		.hps_0_f2h_axi_slave_aruser                                       (mm_interconnect_1_hps_0_f2h_axi_slave_aruser),       //                                                           .aruser
		.hps_0_f2h_axi_slave_arvalid                                      (mm_interconnect_1_hps_0_f2h_axi_slave_arvalid),      //                                                           .arvalid
		.hps_0_f2h_axi_slave_arready                                      (mm_interconnect_1_hps_0_f2h_axi_slave_arready),      //                                                           .arready
		.hps_0_f2h_axi_slave_rid                                          (mm_interconnect_1_hps_0_f2h_axi_slave_rid),          //                                                           .rid
		.hps_0_f2h_axi_slave_rdata                                        (mm_interconnect_1_hps_0_f2h_axi_slave_rdata),        //                                                           .rdata
		.hps_0_f2h_axi_slave_rresp                                        (mm_interconnect_1_hps_0_f2h_axi_slave_rresp),        //                                                           .rresp
		.hps_0_f2h_axi_slave_rlast                                        (mm_interconnect_1_hps_0_f2h_axi_slave_rlast),        //                                                           .rlast
		.hps_0_f2h_axi_slave_rvalid                                       (mm_interconnect_1_hps_0_f2h_axi_slave_rvalid),       //                                                           .rvalid
		.hps_0_f2h_axi_slave_rready                                       (mm_interconnect_1_hps_0_f2h_axi_slave_rready),       //                                                           .rready
		.clk_0_clk_clk                                                    (avalon_clk_clk),                                     //                                                  clk_0_clk.clk
		.avalon_f2h_reset_reset_bridge_in_reset_reset                     (rst_controller_001_reset_out_reset),                 //                     avalon_f2h_reset_reset_bridge_in_reset.reset
		.hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                 // hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.avalon_f2h_avalon_universal_master_0_address                     (avalon_f2h_avalon_universal_master_0_address),       //                       avalon_f2h_avalon_universal_master_0.address
		.avalon_f2h_avalon_universal_master_0_waitrequest                 (avalon_f2h_avalon_universal_master_0_waitrequest),   //                                                           .waitrequest
		.avalon_f2h_avalon_universal_master_0_burstcount                  (avalon_f2h_avalon_universal_master_0_burstcount),    //                                                           .burstcount
		.avalon_f2h_avalon_universal_master_0_byteenable                  (avalon_f2h_avalon_universal_master_0_byteenable),    //                                                           .byteenable
		.avalon_f2h_avalon_universal_master_0_read                        (avalon_f2h_avalon_universal_master_0_read),          //                                                           .read
		.avalon_f2h_avalon_universal_master_0_readdata                    (avalon_f2h_avalon_universal_master_0_readdata),      //                                                           .readdata
		.avalon_f2h_avalon_universal_master_0_readdatavalid               (avalon_f2h_avalon_universal_master_0_readdatavalid), //                                                           .readdatavalid
		.avalon_f2h_avalon_universal_master_0_write                       (avalon_f2h_avalon_universal_master_0_write),         //                                                           .write
		.avalon_f2h_avalon_universal_master_0_writedata                   (avalon_f2h_avalon_universal_master_0_writedata),     //                                                           .writedata
		.avalon_f2h_avalon_universal_master_0_lock                        (avalon_f2h_avalon_universal_master_0_lock),          //                                                           .lock
		.avalon_f2h_avalon_universal_master_0_debugaccess                 (avalon_f2h_avalon_universal_master_0_debugaccess)    //                                                           .debugaccess
	);

	soc_system_mm_interconnect_2 mm_interconnect_2 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                                           //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                                         //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                                          //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                                         //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                                        //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                                         //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                                        //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                                         //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                                        //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                                        //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                                            //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                                          //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                                          //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                                          //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                                         //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                                         //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                                            //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                                          //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                                         //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                                         //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                                           //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                                         //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                                          //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                                         //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                                        //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                                         //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                                        //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                                         //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                                        //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                                        //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                                            //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                                          //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                                          //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                                          //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                                         //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                                         //                                                           .rready
		.clk_1_clk_clk                                                    (avalon_clk_lw_clk),                                                   //                                                  clk_1_clk.clk
		.avalon_h2f_reset_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),                                      //                     avalon_h2f_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                  // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.avalon_h2f_avalon_universal_slave_0_address                      (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_address),       //                        avalon_h2f_avalon_universal_slave_0.address
		.avalon_h2f_avalon_universal_slave_0_write                        (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_write),         //                                                           .write
		.avalon_h2f_avalon_universal_slave_0_read                         (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_read),          //                                                           .read
		.avalon_h2f_avalon_universal_slave_0_readdata                     (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_readdata),      //                                                           .readdata
		.avalon_h2f_avalon_universal_slave_0_writedata                    (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_writedata),     //                                                           .writedata
		.avalon_h2f_avalon_universal_slave_0_burstcount                   (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_burstcount),    //                                                           .burstcount
		.avalon_h2f_avalon_universal_slave_0_byteenable                   (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_byteenable),    //                                                           .byteenable
		.avalon_h2f_avalon_universal_slave_0_readdatavalid                (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_readdatavalid), //                                                           .readdatavalid
		.avalon_h2f_avalon_universal_slave_0_waitrequest                  (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_waitrequest),   //                                                           .waitrequest
		.avalon_h2f_avalon_universal_slave_0_lock                         (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_lock),          //                                                           .lock
		.avalon_h2f_avalon_universal_slave_0_debugaccess                  (mm_interconnect_2_avalon_h2f_avalon_universal_slave_0_debugaccess),   //                                                           .debugaccess
		.h2f_ram_s1_address                                               (mm_interconnect_2_h2f_ram_s1_address),                                //                                                 h2f_ram_s1.address
		.h2f_ram_s1_write                                                 (mm_interconnect_2_h2f_ram_s1_write),                                  //                                                           .write
		.h2f_ram_s1_readdata                                              (mm_interconnect_2_h2f_ram_s1_readdata),                               //                                                           .readdata
		.h2f_ram_s1_writedata                                             (mm_interconnect_2_h2f_ram_s1_writedata),                              //                                                           .writedata
		.h2f_ram_s1_byteenable                                            (mm_interconnect_2_h2f_ram_s1_byteenable),                             //                                                           .byteenable
		.h2f_ram_s1_chipselect                                            (mm_interconnect_2_h2f_ram_s1_chipselect),                             //                                                           .chipselect
		.h2f_ram_s1_clken                                                 (mm_interconnect_2_h2f_ram_s1_clken)                                   //                                                           .clken
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~avalon_reset_lw_reset_n),           // reset_in0.reset
		.clk            (avalon_clk_lw_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~avalon_reset_reset_n),              // reset_in0.reset
		.clk            (avalon_clk_clk),                     //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (avalon_clk_lw_clk),                  //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (avalon_clk_clk),                     //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
